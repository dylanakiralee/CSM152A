`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   03:21:20 03/30/2021
// Design Name:   FPCVT
// Module Name:   /home/ise/CSM152A/Proj1/FPCVT_TB.v
// Project Name:  Proj1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: FPCVT
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module FPCVT_TB;

	// Inputs
	reg [12:0] D;

	// Outputs
	wire S;
	wire [2:0] E;
	wire [4:0] F;

	// Instantiate the Unit Under Test (UUT)
	FPCVT uut (
		.D(D), 
		.S(S), 
		.E(E), 
		.F(F)
	);

	initial begin
		
		D = 13'b0000000000000; // 0
		#10;
		D = 13'b0000000000001; // 1
		#10;
		D = 13'b1111111111111; // -1
		#10;
		D = 13'b1000000000000; //-4096
		#10;
		D = 13'b0111111111111; // 4095
		#10;
		D = 13'b1000000000001; // -4095
		#10;
		D = 13'b0000000000010; // 2
		#10;
		D = 13'b1111111111110; // -2
		#10;
		D = 13'b0000000000011; // 3
		#10;
		D = 13'b1111111111101; // -3
		#10;
		D = 13'b0000000000101; // 5
		#10;
		D = 13'b1111111111011; // -5
		#10;
		D = 13'b0000000001101; // 13
		#10;
		D = 13'b1111111110011; // -13
		#10;
		D = 13'b0000000011001; // 25
		#10;
		D = 13'b1111111100111; // -25
		#10;
		D = 13'b0000000111111; // 63
		#10;
		D = 13'b1111111000001; // -63
		#10;
		D = 13'b0000001011101; // 93
		#10;
		D = 13'b1111110100011; // -93
		#10;
		D = 13'b0000010011001; // 153
		#10;
		D = 13'b1111101100111; // -153
		#10;
		D = 13'b0000101011001; // 345
		#10;
		D = 13'b1111010100111; // -345
		#10;
		D = 13'b0001101011101; // 861
		#10;
		D = 13'b1110010100011; // -861
		#10;
		D = 13'b0010101011101; // 1373
		#10;
		D = 13'b1101010100011; // -1373
		#10;
		D = 13'b0110101011100; // 3420
		#10;
		D = 13'b1001010100100; // -3420
		#10;
	end
      
endmodule

